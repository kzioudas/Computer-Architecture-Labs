-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Wed Oct 31 13:26:26 2018"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY regCmp IS 
	PORT
	(
		true_wren :  IN  STD_LOGIC;
		ra :  IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		wa :  IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		bypass :  OUT  STD_LOGIC
	);
END regCmp;

ARCHITECTURE bdf_type OF regCmp IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_2 <= NOT(ra(4) XOR wa(4));


SYNTHESIZED_WIRE_3 <= NOT(ra(3) XOR wa(3));


SYNTHESIZED_WIRE_0 <= NOT(ra(1) XOR wa(1));


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_0 AND SYNTHESIZED_WIRE_1 AND true_wren;


SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_2 AND SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_4;


bypass <= SYNTHESIZED_WIRE_5 AND SYNTHESIZED_WIRE_6;


SYNTHESIZED_WIRE_4 <= NOT(ra(2) XOR wa(2));


SYNTHESIZED_WIRE_1 <= NOT(ra(0) XOR wa(0));


END bdf_type;